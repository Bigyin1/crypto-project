
module crypto(input logic clk_i);


endmodule
